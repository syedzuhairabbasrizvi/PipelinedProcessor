`timescale 1ns / 1ps
module instruction_parser(
    input [31:0] instruction,
    output [6:0] opcode,
    output [4:0] rd,
    output [2:0] funct3,
    output [4:0] rs1,
    output [4:0] rs2,
    output [6:0] funct7
);
//simple: just slice instruction accordingly as per R format
/*
assign opcode = instruction[6:0];
assign rd = instruction[11:7];
assign funct3 = instruction[14:12];
assign rs1 = instruction[19:15];
assign rs2 = instruction[24:20];
assign funct7 = instruction[31:25];
*/
// Extracting opcode
assign opcode = instruction[6:0];

// Determining instruction format using opcode
assign {rd, funct3, rs1, rs2, funct7} = (opcode == 7'b0110011) ? // R format
                                        {instruction[11:7], instruction[14:12], instruction[19:15], instruction[24:20], instruction[31:25]} :
                                        (opcode == 7'b0000011 | opcode == 7'b0010011) ? // I format
                                        {instruction[11:7], instruction[14:12], instruction[19:15], 5'b0, 7'b0} :
                                        // Assuming opcode for S format is 7'b0100011
                                        {5'b0, instruction[14:12], instruction[19:15], instruction[24:20], 7'b0};

endmodule


